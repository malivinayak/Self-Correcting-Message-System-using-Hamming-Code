module vinayak_inverter(output Y, input A);
    not (Y, A);
endmodule